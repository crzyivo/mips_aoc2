----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:38:18 05/15/2014 
-- Design Name: 
-- Module Name:    UC_slave - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: la UC incluye un contador de 2 bits para llevar la cuenta de las transferencias de bloque y una m�quina de estados
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity UC_MC is
    Port ( 	clk : in  STD_LOGIC;
			reset : in  STD_LOGIC;
			RE : in  STD_LOGIC; --RE y WE son las ordenes del MIPs
			WE : in  STD_LOGIC;
			hit : in  STD_LOGIC; --se activa si hay acierto
			bus_TRDY : in  STD_LOGIC; --indica que la memoria no puede realizar la operaci�n solicitada en este ciclo
			Bus_DevSel: in  STD_LOGIC; --indica que la memoria ha reconocido que la direcci�n est� dentro de su rango
			MC_RE : out  STD_LOGIC; --RE y WE de la MC
            MC_WE : out  STD_LOGIC;
            MC_bus_Rd_Wr : out  STD_LOGIC; --1 para escritura en Memoria y 0 para lectura
            MC_tags_WE : out  STD_LOGIC; -- para escribir la etiqueta en la memoria de etiquetas
            palabra : out  STD_LOGIC_VECTOR (1 downto 0);--indica la palabra actual dentro de una transferencia de bloque (1�, 2�...)
            mux_origen: out STD_LOGIC; -- Se utiliza para elegir si el origen de la direcci�n y el dato es el Mips (cuando vale 0) o la UC y el bus (cuando vale 1)
            ready : out  STD_LOGIC; -- indica si podemos procesar la orden actual del MIPS en este ciclo. En caso contrario habr� que detener el MIPs
            block_addr : out  STD_LOGIC; -- indica si la direcci�n a enviar es la de bloque (rm) o la de palabra (w)
			MC_send_addr : out  STD_LOGIC; --ordena que se env�en la direcci�n y las se�ales de control al bus
            MC_send_data : out  STD_LOGIC; --ordena que se env�en los datos
            Frame : out  STD_LOGIC; --indica que la operaci�n no ha terminado
			Replace_block	: out  STD_LOGIC; -- indica que se ha reemplazado un bloque
			inc_rm : out STD_LOGIC; -- indica que ha habido un fallo de lectura
			inc_wm : out STD_LOGIC; -- indica que ha habido un fallo de escritura
			inc_wh : out STD_LOGIC -- indica que ha habido un acierto de escritura
           );
end UC_MC;

architecture Behavioral of UC_MC is


component counter_2bits is
		    Port ( clk : in  STD_LOGIC;
		           reset : in  STD_LOGIC;
		           count_enable : in  STD_LOGIC;
		           count : out  STD_LOGIC_VECTOR (1 downto 0)
					  );
end component;		           
-------------------------------------------------------------------------------------------------
-- poner en el siguiente type el nombre de vuestros estados
type state_type is (Inicio, MD_write,MD_write_rdy,MD_read_rdy,MD_read,Cooldown); 
signal state, next_state : state_type; 
signal last_word: STD_LOGIC; --se activa cuando se est� pidiendo la �ltima palabra de un bloque
signal count_enable: STD_LOGIC; -- se activa si se ha recibido una palabra de un bloque para que se incremente el contador de palabras
signal palabra_UC : STD_LOGIC_VECTOR (1 downto 0);
begin
 
 
--el contador nos dice cuantas palabras hemos recibido. Se usa para saber cuando se termina la transferencia del bloque y para direccionar la palabra en la que se escribe el dato leido del bus en la MC
word_counter: counter_2bits port map (clk, reset, count_enable, palabra_UC); --indica la palabra actual dentro de una transferencia de bloque (1�, 2�...)

last_word <= '1' when palabra_UC="11" else '0';--se activa cuando estamos pidiendo la �ltima palabra

palabra <= palabra_UC;

   SYNC_PROC: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (reset = '1') then
            state <= Inicio;
         else
            state <= next_state;
         end if;        
      end if;
   end process;
 

   -- Poned aqu� el c�digo de vuestra m�quina de estados
   OUTPUT_DECODE: process (state, hit, last_word, bus_TRDY, RE, WE, Bus_DevSel)
   begin
		-- Se comienza dando los valores por defecto, si no se asigna otro valor en un estado valdr�n lo que se asigna aqu�
		-- As� no hay que asignar valor a todas las se�ales en cada caso
		MC_WE <= '0';
		MC_bus_Rd_Wr <= '0';
		MC_tags_WE <= '0';
        MC_RE <= RE;
        ready <= '0';
        mux_origen <= '0';
        MC_send_addr <= '0';
        MC_send_data <= '0';
        next_state <= state;  
		count_enable <= '0';
		Frame <= '0';
		Replace_block <= '0';	
		block_addr <= '0';
		inc_rm <= '0';
		inc_wm <= '0';
		inc_wh <= '0';
			
        -- Estado Inicio          
        if (state = Inicio and RE= '0' and WE= '0') then -- si no piden nada no hacemos nada
				next_state <= Inicio;
				ready <= '1';

		elsif (state = Inicio and WE='1' and hit='0') then --Tenemos fallo en escritura, escribimos directamente en MD
					ready <= '0';
					Frame <='1';
					next_state <= MD_write_rdy;
					MC_bus_Rd_Wr <= '1';
					MC_send_addr <='1';
					inc_wm <='1';

		elsif (state=Inicio and RE= '1' and hit='0') then --Tenemos fallo en lectura, paramos y pedimos bloque a MD
					ready <='0';
					MC_send_addr <='1';
					next_state <= MD_read_rdy;
					inc_rm <='1';
					block_addr <='1';

		elsif (state=Inicio and hit='1') then --Tenemos acierto
				ready <= '1';
				next_state <= Inicio; --Si resulta acierto, pero ha sido casualidad, no hacemos nada mas
				if(RE='1') then
					MC_RE <= '1'; --Si era acierto en lectura, leemos de cache y vale
				end if;
				if(WE='1') then --Si es acierto de escritura, escribimos en cache y paramos hasta haber realizado la escritura en MD
					ready <= '0';
					Frame <='1';
					next_state <= MD_write_rdy;
					MC_WE<= '1';
					MC_bus_Rd_Wr <= '1';
					MC_send_addr <='1';
					inc_wh <='1';
				end if;

--------------------------------------------Escrituras: MD_write_rdy y MD_write------------------------------------------------------------------------				
		elsif (state=MD_write_rdy and Bus_DevSel='0') then --Se realiza una escritura en MD, pero aun no esta listo MD
				Frame <='1';
				next_state <= MD_write_rdy;
				MC_bus_Rd_Wr <= '1';
				MC_send_addr <='1';
		elsif (state=MD_write_rdy and Bus_DevSel='1') then --Se realiza escritura y se reconoze la direccion, procedemos a enviar dato
				Frame <='1';
				next_state <= MD_write;
				MC_bus_Rd_Wr <='1';
				MC_send_data <= '1';

		elsif (state=MD_write and bus_TRDY='1') then --Se realiza la escritura en MD, volvemos a Inicio y dejamos continuar a MIPS
				next_state <=Cooldown;
				Frame <= '1';
				MC_bus_Rd_Wr <='1';
				MC_send_data <= '1';
		elsif (state=MD_write and bus_TRDY='0') then --MD no esta lista para escribir, mantenemos el dato en el bus
				next_state<= MD_write;
				Frame <='1';
				MC_bus_Rd_Wr <='1';
				MC_send_data <= '1';

		--------------------------------------------Fallo Lectura: MD_read_rdy y MD_read------------------------------------------------------------------------
		elsif (state=MD_read_rdy and Bus_DevSel='0') then --MD no esta lista para mandar el bloque
				next_state <= MD_read_rdy;
				Frame <= '1';
				MC_send_addr <= '1';
				block_addr <='1';
		elsif(state=MD_read_rdy and Bus_DevSel='1') then --MD lista para mandar el bloque
				next_state <= MD_read;
				Frame <='1';

		elsif (state=MD_read and bus_TRDY='0') then --Retardo en el envio de la palabra
				Frame <='1';
				next_state <=MD_read;
		elsif (state=MD_read and bus_TRDY='1') then --Se envia la palabra desde MD, si es la primera escribimos el TAG
				Frame <='1';
				next_state <=MD_read;
				MC_WE <= '1';
				mux_origen <='1';
				count_enable <='1';
				if(palabra_UC="00") then --Primera palabra recibida, actualizo tags
					MC_tags_WE <='1';
				end if;
				if(last_word='1') then --Fin de recepcion de bloque
					next_state <= Cooldown;
					Replace_block <='1';
				end if;
--------------------------------------------CoolDown------------------------------------------------------------------------				
		elsif (state=Cooldown) then --Ciclo extra para mantener Frame a 0 y no confundir a MD_cont
				next_state<=Inicio;
				Frame <='0';
		end if;
   end process;
 
   
end Behavioral;